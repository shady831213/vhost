 `ifndef __MAILBOX_SVH__
 `define __MAILBOX_SVH__
 `ifndef MB_PTR
 `define MB_PTR longint unsigned
 `endif
`ifndef SV_CALL_MAX_ARGS
 `define SV_CALL_MAX_ARGS 16
`endif
`endif
