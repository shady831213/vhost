`ifndef __MAILBOX_IF_SV__
`define __MAILBOX_IF_SV__
interface MailboxIf();
   bit clk;
   bit reset;
endinterface
`endif
